library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

ENTITY dds_gen_yt IS
  GENERIC (
    addr_width : integer := 8;      -- 2^8 = 256 LUT-Schritte
    data_width : integer := 16;
    clk_freq   : integer := 48000;  -- Hz
    out_freq   : integer := 1319    -- Hz
  );
  PORT (
    clk, reset : in std_logic;
    data_a     : out std_logic_vector(data_width-1 downto 0)
  );
END dds_gen_yt;

ARCHITECTURE arch OF dds_gen_yt IS

  constant PHASE_WIDTH : integer := 24;  -- DDS: Großer Phase-Accu!

  type LUT_TYPE is array (0 to 255) of integer;
  constant LUT : LUT_TYPE := (
  0,
184,369,554,738,923,1107,1291,1476,1659,1843,2026,2209,2392,2574,2756,2937,3118,3299,3479,3658,
3837,4015,4193,4370,4547,4723,4898,5072,5245,5418,5590,5761,5931,6101,6269,6436,6603,6768,6933,7096,
7258,7419,7579,7738,7896,8052,8208,8362,8515,8666,8816,8965,9113,9259,9403,9547,9688,9829,9968,10105,
10241,10375,10508,10639,10768,10896,11022,11147,11269,11391,11510,11628,11743,11857,11970,12080,12189,12296,12401,12504,
12605,12704,12801,12896,12990,13081,13171,13258,13344,13427,13508,13588,13665,13740,13813,13884,13953,14020,14084,14147,
14207,14265,14321,14375,14427,14476,14524,14569,14612,14652,14691,14727,14761,14793,14822,14849,14874,14897,14917,14936,
14951,14965,14976,14986,14992,14997,14999,14999,14997,14992,14986,14976,14965,14951,14936,14917,14897,14874,14849,14822,
14793,14761,14727,14691,14652,14612,14569,14524,14476,14427,14375,14321,14265,14207,14147,14084,14020,13953,13884,13813,
13740,13665,13588,13508,13427,13344,13258,13171,13081,12990,12896,12801,12704,12605,12504,12401,12296,12189,12080,11970,
11857,11743,11628,11510,11391,11269,11147,11022,10896,10768,10639,10508,10375,10241,10105,9968,9829,9688,9547,9403,
9259,9113,8965,8816,8666,8515,8362,8208,8052,7896,7738,7579,7419,7258,7096,6933,6768,6603,6436,6269,
6101,5931,5761,5590,5418,5245,5072,4898,4723,4547,4370,4193,4015,3837,3658,3479,3299,3118,2937,2756,
2574,2392,2209,2026,1843,1659,1476,1291,1107,923,738,554,369,184,0
  );

  constant PHASE_INC : unsigned(PHASE_WIDTH-1 downto 0) :=
    to_unsigned(integer(2**PHASE_WIDTH * out_freq / (clk_freq*10)), PHASE_WIDTH);

  signal phase_acc : unsigned(PHASE_WIDTH-1 downto 0) := (others => '0');
  signal lut_addr  : integer range 0 to 255 := 0;

BEGIN

  data_a <= std_logic_vector(to_unsigned(LUT(lut_addr), data_width));

  PROCESS(clk, reset)
  BEGIN
    IF reset = '1' THEN
      phase_acc <= (others => '0');
    ELSIF rising_edge(clk) THEN
      phase_acc <= phase_acc + PHASE_INC;

      lut_addr <= to_integer(phase_acc(PHASE_WIDTH-1 downto PHASE_WIDTH-addr_width));
    END IF;
  END PROCESS;

END arch;
